// megafunction wizard: %ALTFP_INV%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTFP_INV 

// ============================================================
// File Name: invert.v
// Megafunction Name(s):
// 			ALTFP_INV
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.1.0 Build 590 10/25/2017 SJ Lite Edition
// ************************************************************

//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

module invert (
	clock,
	data,
	result)/* synthesis synthesis_clearbox = 1 */;

	input	  clock;
	input	[31:0]  data;
	output	[31:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_inv"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "20"
// Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
// Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
// Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
// Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
// Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
// Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL invert.cmp TRUE TRUE
// Retrieval info: LIB_FILE: lpm
